library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity buffered_vga is
    port (
        a: in integer
    );
end entity buffered_vga;

architecture behav of buffered_vga is
    
begin
    
end architecture behav;